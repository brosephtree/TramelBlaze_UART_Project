`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/01/2020 05:13:35 PM
// Design Name: 
// Module Name: led_module
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module led_module(
    input clock,
    input reset,
    input D,
    input LD,
    output [15:0] led
    );
    
    parameter CLK_FREQ = 100 * 10**6;           //clock at 100 MHz
    
    
    
    
    
endmodule
